


parameter ADD = 3'b000;
parameter SUB = 3'b001;
parameter SLL = 3'b010;
parameter SLT = 3'b011;
parameter SRL = 3'b100;
parameter XOR_= 3'b101;
parameter OR_ = 3'b110;
parameter AND_= 3'b111;

parameter LW = 7'b0000011;
parameter SW = 7'b0100011;
parameter R_type = 7'b0110011;
parameter I_type = 7'b0010011;
parameter JAL = 7'b1101111;
parameter BEQ = 7'b1100011;
